module mul(input logic [7:0] a, b, output logic [7:0] product);
    assign product = a*b;
endmodule