module none();
endmodule