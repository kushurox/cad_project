module mul(input logic [3:0] a, b, output logic [3:0] product);
    assign product = a*b;
endmodule